module routes

import structs { App }

pub struct AliasApp {
	App
}
