module api

import structs { App }

pub struct Api {
	App
}
