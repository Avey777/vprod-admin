module tenant_api

import internal.structs { App }

pub struct Api {
	App
}
