module tenant_menu

import internal.structs { App }

pub struct Menu {
	App
}
