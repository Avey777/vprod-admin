module fms_api

import structs { App }

type HandlerApp = App
