module handler

import log
import admin { Admin }

pub fn register_routes(mut app App) {
	mut admin_app := &Admin{}

	app.register_controller[Admin, Context]('/admin', mut admin_app) or { log.error('${err}') }
}

pub fn before_request(mut ctx Context) bool {
	// $if trace_before_request ? {
	log.info('[veb] before_request: ${ctx.req.method} ${ctx.req.url}')
	// }
	return true
}
