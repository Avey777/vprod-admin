// role_permission | authority | 角色权限分配和获取

module role_permission

import structs { App }

pub struct RolePermission {
	App
}
