module token

import internal.structs { App }

pub struct Token {
	App
}
