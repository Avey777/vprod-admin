module authentication

import internal.structs { App }

pub struct Authentication {
	App
}
