module token

import structs { App }

pub struct Token {
	App
}
