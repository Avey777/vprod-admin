module base_api

import internal.structs { App }

type HandlerApp = App
