module route

import structs { App }

pub struct AliasApp {
	App
}
