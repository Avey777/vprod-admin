module oauthprovider

import structs { App }

pub struct OauthProvider {
	App
}
