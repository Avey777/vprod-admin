module tasklog

// import (
// 	"context"

// 	"github.com/suyuan32/simple-admin-common/i18n"
// 	"github.com/zeromicro/go-zero/core/errorx"

// 	"github.com/suyuan32/simple-admin-job/types/job"

// 	"github.com/suyuan32/simple-admin-core/api/internal/svc"
// 	"github.com/suyuan32/simple-admin-core/api/internal/types"

// 	"github.com/zeromicro/go-zero/core/logx"
// )

// type CreateTaskLogLogic struct {
// 	logx.Logger
// 	ctx    context.Context
// 	svcCtx *svc.ServiceContext
// }

// func NewCreateTaskLogLogic(ctx context.Context, svcCtx *svc.ServiceContext) *CreateTaskLogLogic {
// 	return &CreateTaskLogLogic{
// 		Logger: logx.WithContext(ctx),
// 		ctx:    ctx,
// 		svcCtx: svcCtx,
// 	}
// }

// func (l *CreateTaskLogLogic) CreateTaskLog(req *types.TaskLogInfo) (resp *types.BaseMsgResp, err error) {
// 	if !l.svcCtx.Config.JobRpc.Enabled {
// 		return nil, errorx.NewCodeUnavailableError(i18n.ServiceUnavailable)
// 	}
// 	data, err := l.svcCtx.JobRpc.CreateTaskLog(l.ctx,
// 		&job.TaskLogInfo{
// 			StartedAt:  req.StartedAt,
// 			FinishedAt: req.FinishedAt,
// 			Result:     req.Result,
// 		})
// 	if err != nil {
// 		return nil, err
// 	}
// 	return &types.BaseMsgResp{Msg: l.svcCtx.Trans.Trans(l.ctx, data.Msg)}, nil
// }
