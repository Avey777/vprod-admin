module api

import veb
import log
import time
import orm
import x.json2
import internal.structs.schema_sys
import common.api
import internal.structs { Context }

@['/list'; post]
fn (app &Api) api_list(mut ctx Context) veb.Result {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')
	// log.debug('ctx.req.data type: ${typeof(ctx.req.data).name}')

	req := json2.raw_decode(ctx.req.data) or { return ctx.json(api.json_error_400(err.msg())) }
	mut result := api_list_resp(mut ctx, req) or { return ctx.json(api.json_error_500(err.msg())) }

	return ctx.json(api.json_success_200(result))
}

fn api_list_resp(mut ctx Context, req json2.Any) !map[string]Any {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	page := req.as_map()['page'] or { 1 }.int()
	page_size := req.as_map()['page_size'] or { 10 }.int()
	path := req.as_map()['path'] or { '' }.str()
	api_group := req.as_map()['api_group'] or { '' }.str()
	service_name := req.as_map()['service_name'] or { '' }.str()
	method := req.as_map()['method'] or { '' }.str()
	is_required := req.as_map()['is_required'] or { 100 }.u8()

	db, conn := ctx.dbpool.acquire() or { return error('Failed to acquire connection: ${err}') }
	defer {
		ctx.dbpool.release(conn) or {
			log.warn('Failed to release connection ${@LOCATION}: ${err}')
		}
	}

	mut sys_api := orm.new_query[schema_sys.SysApi](db)
	// 总页数查询 - 分页偏移量构造
	mut count := sql db {
		select count from schema_sys.SysUser
	}!
	offset_num := (page - 1) * page_size
	//*>>>*/
	mut query := sys_api.select()!
	if path != '' {
		query = query.where('path = ?', path)!
	}
	if api_group != '' {
		query = query.where('api_group = ?', api_group)!
	}
	if service_name != '' {
		query = query.where('service_name = ?', service_name)!
	}
	if is_required !in [0, 1] {
		query = query.where('is_required = ?', is_required)!
	}
	if method != '' {
		query = query.where('method = ?', method)!
	}

	result := query.limit(page_size)!.offset(offset_num)!.query()!
	//*<<<*/
	mut datalist := []map[string]Any{} // map空数组初始化
	for row in result {
		mut data := map[string]Any{} // map初始化
		data['id'] = row.id //主键ID
		data['path'] = row.path
		data['description'] = row.description or { '' }
		data['api_group'] = row.api_group
		data['method'] = row.method
		data['is_required'] = int(row.is_required)
		data['service_name'] = row.service_name

		data['created_at'] = row.created_at.format_ss()
		data['updated_at'] = row.updated_at.format_ss()
		data['deleted_at'] = row.deleted_at or { time.Time{} }.format_ss()

		datalist << data //追加data到maplist 数组
	}

	mut result_data := map[string]Any{}
	result_data['total'] = count
	result_data['data'] = datalist

	return result_data
}
