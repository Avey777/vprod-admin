module config

// import internal.config

// fn test_set_web_port() {
// 	web_port := config.set_web_port()
// 	assert typeof(web_port).name == 'int'
// 	assert web_port > 1000 && web_port < 65535
// }
