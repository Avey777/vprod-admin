module user

import internal.structs { App }

pub struct User {
	App
}
