module role

import structs { App }

pub struct Role {
	App
}
