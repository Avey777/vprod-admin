module department

import veb
import log
import orm
import x.json2
import internal.config { db_mysql }
import internal.structs.schema
import internal.structs { Context, json_error, json_success }

// Delete department | 删除department
@['/delete_department'; post]
fn (app &Department) delete_department(mut ctx Context) veb.Result {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	req := json2.raw_decode(ctx.req.data) or { return ctx.json(json_error(502, '${err}')) }
	mut result := delete_department_resp(req) or { return ctx.json(json_error(503, '${err}')) }

	return ctx.json(json_success('success', result))
}

fn delete_department_resp(req json2.Any) !map[string]Any {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	mut db := db_mysql()
	defer { db.close() }

	department_id := req.as_map()['id'] or { '' }.str()

	mut sys_department := orm.new_query[schema.SysDepartment](db)
	sys_department.delete()!.where('id = ?', department_id)!.update()!
	// sys_department.set('del_flag = ?', 1)!.where('id = ?', department_id)!.update()!

	return map[string]Any{}
}
