module api

import veb
// import pool

pub struct Context {
	veb.Context
}
