module project

import structs { App }

pub struct Project {
	App
}
