module menu

import internal.structs { App }

pub struct Menu {
	App
}
