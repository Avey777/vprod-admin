// role_permission | 角色权限分配和获取

module authority

import internal.structs { App }

pub struct RolePermission {
	App
}
