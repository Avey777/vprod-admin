module db_api

import structs { App }

pub struct Base {
	App
}
