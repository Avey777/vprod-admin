module routes

import internal.structs { App }

pub struct AliasApp {
	App
}
