module api

import internal.structs { App }

pub struct Api {
	App
}
