module role

import internal.structs { App }

pub struct Role {
	App
}
