module i18n

import time
import os
import log
import x.json2 as json

// ------------------------- I18n -------------------------
@[heap]
pub struct I18nStore {
pub:
	default_lang string
	dir          string
pub mut:
	translations   map[string]map[string]string
	lang_cache     map[string]string
	mod_times      map[string]int
	last_check     i64
	check_interval i64 = 2000 // 毫秒
}

// 创建 I18nStore
pub fn new_i18n(dir string, default_lang string) !&I18nStore {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	mut s := &I18nStore{
		dir:          dir
		default_lang: default_lang
		translations: map[string]map[string]string{}
		lang_cache:   map[string]string{}
		mod_times:    map[string]int{}
		last_check:   0
	}
	load_translations(mut s)!
	return s
}

// ------------------------- 动态加载 + JSON 校验 + 日志 -------------------------
pub fn maybe_reload(mut s I18nStore) {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	now := time.now().unix()
	if now - s.last_check < s.check_interval / 1000 {
		return
	}
	s.last_check = now
	load_translations(mut s) or { eprintln('i18n load failed: ${err}') }
}

pub fn load_translations(mut s I18nStore) ! {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	if !os.exists(s.dir) {
		return
	}
	for file in os.ls(s.dir)! {
		if !file.ends_with('.json') {
			continue
		}
		full_path := os.join_path(s.dir, file)
		mod_time := int(os.file_last_mod_unix(full_path))

		if file in s.mod_times && s.mod_times[file] == mod_time {
			continue
		}

		content := os.read_file(full_path)!

		// JSON 解码，失败则跳过文件
		data := json.decode[map[string]json.Any](content) or {
			eprintln('i18n load failed for ${file}: ${err}')
			continue
		}

		lang := file.replace('.json', '')

		mut is_new := false
		if lang !in s.translations {
			s.translations[lang] = map[string]string{}
			is_new = true
		}

		flat := flatten_map(data, '')
		for k, v in flat {
			s.translations[lang][k] = v
		}

		s.mod_times[file] = mod_time

		// 打印加载日志
		println('i18n loaded: ${lang}, keys: ${s.translations[lang].len}, new: ${is_new}')
	}
}

// 查询翻译，支持 fallback
pub fn (s &I18nStore) t(lang string, key string) string {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	selected := if lang in s.translations.keys() { lang } else { s.default_lang }

	if key in s.translations[selected] {
		return s.translations[selected][key]
	}
	if key in s.translations[s.default_lang] {
		return s.translations[s.default_lang][key]
	}
	return key
}

// 展平成点号路径
fn flatten_map(data map[string]json.Any, prefix string) map[string]string {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	mut result := map[string]string{}
	for k, v in data {
		full_key := if prefix == '' { k } else { '${prefix}.${k}' }
		match v {
			string {
				result[full_key] = v
			}
			map[string]json.Any {
				sub := flatten_map(v, full_key)
				for sk, sv in sub {
					result[sk] = sv
				}
			}
			else {}
		}
	}
	return result
}
