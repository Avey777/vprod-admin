module routes

import internal.structs { App }

pub type AliasApp = App
