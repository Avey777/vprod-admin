module sys_admin

import internal.structs { App }

pub struct Admin {
	App
}
