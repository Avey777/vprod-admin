module structt

import veb

pub struct Context {
	veb.Context
}
