module application

import internal.structs { App }

pub struct Application {
	App
}
