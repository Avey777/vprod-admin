module oauthprovider

import internal.structs { App }

pub struct OauthProvider {
	App
}
