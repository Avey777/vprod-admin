module authentication

// import (
// 	"context"

// 	"github.com/suyuan32/simple-admin-common/config"
// 	"github.com/suyuan32/simple-admin-common/enum/errorcode"
// 	"github.com/suyuan32/simple-admin-common/orm/ent/entctx/datapermctx"
// 	"github.com/suyuan32/simple-admin-common/orm/ent/entenum"
// 	"github.com/suyuan32/simple-admin-common/utils/pointy"
// 	"github.com/zeromicro/go-zero/core/errorx"

// 	"github.com/suyuan32/simple-admin-core/api/internal/svc"
// 	"github.com/suyuan32/simple-admin-core/api/internal/types"
// 	"github.com/suyuan32/simple-admin-core/rpc/types/core"

// 	"github.com/zeromicro/go-zero/core/logx"
// )

// type RegisterLogic struct {
// 	logx.Logger
// 	ctx    context.Context
// 	svcCtx *svc.ServiceContext
// }

// func NewRegisterLogic(ctx context.Context, svcCtx *svc.ServiceContext) *RegisterLogic {
// 	return &RegisterLogic{
// 		Logger: logx.WithContext(ctx),
// 		ctx:    ctx,
// 		svcCtx: svcCtx,
// 	}
// }

// func (l *RegisterLogic) Register(req *types.RegisterReq) (resp *types.BaseMsgResp, err error) {
// 	if l.svcCtx.Config.ProjectConf.RegisterVerify != "captcha" {
// 		return nil, errorx.NewCodeAbortedError("login.registerTypeForbidden")
// 	}

// 	if ok := l.svcCtx.Captcha.Verify(config.RedisCaptchaPrefix+req.CaptchaId, req.Captcha, true); ok {
// 		l.ctx = datapermctx.WithScopeContext(l.ctx, entenum.DataPermAllStr)

// 		_, err := l.svcCtx.CoreRpc.CreateUser(l.ctx,
// 			&core.UserInfo{
// 				Username:     &req.Username,
// 				Password:     &req.Password,
// 				Email:        &req.Email,
// 				Nickname:     &req.Username,
// 				Status:       pointy.GetPointer(uint32(1)),
// 				HomePath:     pointy.GetPointer("/dashboard"),
// 				RoleIds:      []uint64{l.svcCtx.Config.ProjectConf.DefaultRoleId},
// 				DepartmentId: pointy.GetPointer(l.svcCtx.Config.ProjectConf.DefaultDepartmentId),
// 				PositionIds:  []uint64{l.svcCtx.Config.ProjectConf.DefaultPositionId},
// 			})
// 		if err != nil {
// 			return nil, err
// 		}

// 		resp = &types.BaseMsgResp{
// 			Msg: l.svcCtx.Trans.Trans(l.ctx, "login.signupSuccessTitle"),
// 		}
// 		return resp, nil
// 	} else {
// 		return nil, errorx.NewCodeError(errorcode.InvalidArgument,
// 			l.svcCtx.Trans.Trans(l.ctx, "login.wrongCaptcha"))
// 	}
// }
