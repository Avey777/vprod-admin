module user

import structs { App }

pub struct User {
	App
}
