module application

import structs { App }

pub struct Application {
	App
}
