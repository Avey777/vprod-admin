module authentication

import structs { App }

pub struct Authentication {
	App
}
