module schema
