module mq
