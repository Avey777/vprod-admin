module oauthprovider

import internal.structs { App }

pub struct Oauthprovider {
	App
}
