module db_api

import internal.structs { App }

pub struct Base {
	App
}
