module authentication

import time
import internal.structs { App }

pub struct Authentication {
	App
}
