module handler

import internal.structs { App }

pub type HandlerApp = App
