module main

pub fn banner() {
	cyan := '\x1b[38;5;51m'
	reset := '\x1b[0m'

	println(
		r'
██╗   ██╗    █████╗ ██████╗ ███╗   ███╗██╗███╗   ██╗
██║   ██║   ██╔══██╗██╔══██╗████╗ ████║██║████╗  ██║
██║   ██║   ███████║██║  ██║██╔████╔██║██║██╔██╗ ██║
╚██╗ ██╔╝   ██╔══██║██║  ██║██║╚██╔╝██║██║██║╚██╗██║
 ╚████╔╝    ██║  ██║██████╔╝██║ ╚═╝ ██║██║██║ ╚████║
  ╚═══╝     ╚═╝  ╚═╝╚═════╝ ╚═╝     ╚═╝╚═╝╚═╝  ╚═══╝
' +
		reset)

	println(cyan + ':: v-admin ::    Professional Admin Dashboard (v0.5.0)' + reset)
}
