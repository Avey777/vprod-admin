module logic

import veb

struct Context {
	veb.Context
}

pub struct Admin {}
