module dictionarydetail

import veb
import log
import orm
import x.json2

import internal.structs.schema_sys
import common.api { json_success, json_error }
import internal.structs { Context }

// Delete dictionarydetail | 删除dictionarydetail
@['/delete_dictionarydetail'; post]
fn (app &DictionaryDetail) delete_dictionarydetail(mut ctx Context) veb.Result {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	req := json2.raw_decode(ctx.req.data) or { return ctx.json(api.json_error_400(err.msg())) }
	mut result := delete_dictionarydetail_resp(mut ctx, req) or {
		return ctx.json(api.json_error_500(err.msg()) )
	}

	return ctx.json(api.json_success_200(result) )
}

fn delete_dictionarydetail_resp(mut ctx Context,req json2.Any) !map[string]Any {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	db, conn := ctx.dbpool.acquire() or { return error('Failed to acquire connection: ${err}') }
	defer {
		ctx.dbpool.release(conn) or {
			log.warn('Failed to release connection ${@LOCATION}: ${err}')
		}
	}

	dictionarydetail_id := req.as_map()['id'] or { '' }.str()

	mut sys_dictionarydetail := orm.new_query[schema_sys.SysDictionaryDetail](db)
	sys_dictionarydetail.delete()!.where('id = ?', dictionarydetail_id)!.update()!
	// sys_dictionarydetail.set('del_flag = ?', 1)!.where('id = ?', dictionarydetail_id)!.update()!

	return map[string]Any{}
}
