module base_api

import structs { App }

type HandlerApp = App
