module admin

import structs { App }

pub struct Admin {
	App
}
