module schema

// import time

// // 任务日志表
// @[table: 'task_logs']
// pub struct TaskLog {
// pub:
// 	id                          u64              @[comment: "ID"]
// 	started_at                  time.Time        @[immutable; default: ''; comment: "Task Started Time | 任务启动时间"]
// 	finished_at                 ?time.Time       @[comment: "Task Finished Time | 任务完成时间"]
// 	result                      u8               @[comment: "The Task Process Result | 任务执行结果"]
// }
