module menu

import structs { App }

pub struct Menu {
	App
}
