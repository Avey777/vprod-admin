module project

import internal.structs { App }

pub struct Project {
	App
}
