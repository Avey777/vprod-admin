module user

import internal.structs { App }

pub struct Api {
	App
}
