module sys_admin

import structs { App }

pub struct Admin {
	App
}
