module schema

// import time
// import rand

// // 任务表
// @[table: 'tasks']
// pub struct Task {
// pub:
//   id                          uuid        @[immutable; default: ''] // UUID

// 	name                        string           @[comment: "Task Name | 任务名称"]
// 	task_group                  string           @[comment: "Task Group | 任务分组"]
// 	cron_expression             string           @[comment: "Cron expression | 定时任务表达式"]
// 	pattern                     string           @[comment: "Cron Pattern | 任务的模式 （用于区分和确定要执行的任务）"]
// 	payload                     string           @[comment: "The data used in cron (JSON string) | 任务需要的数据(JSON 字符串)"]
// }
