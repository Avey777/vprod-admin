module role_permission

import internal.structs { App }

pub struct RolePermission {
	App
}
