module tenant

import internal.structs { App }

pub struct Tenant {
	App
}
