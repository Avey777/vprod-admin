module role

import veb
import log
import orm
import x.json2 as json
import structs.schema_core { CoreRole }
import common.api
import structs { Context }

// ----------------- Handler 层 -----------------
@['/tenant_role/delete'; post]
pub fn delete_role_handler(app &Role, mut ctx Context) veb.Result {
	log.debug('${@METHOD}  ${@MOD}.${@FILE_LINE}')

	req := json.decode[DeleteTenantRoleReq](ctx.req.data) or {
		return ctx.json(api.json_error_400(err.msg()))
	}

	result := delete_role_usecase(mut ctx, req) or {
		return ctx.json(api.json_error_500('Internal Server Error: ${err}'))
	}

	return ctx.json(api.json_success_200(result))
}

// ----------------- Application Service | Usecase 层 -----------------
pub fn delete_role_usecase(mut ctx Context, req DeleteTenantRoleReq) !DeleteTenantRoleResp {
	// 参数校验
	delete_role_domain(req)!

	// 执行删除
	return delete_role_repo(mut ctx, req)
}

// ----------------- Domain 层 -----------------
fn delete_role_domain(req DeleteTenantRoleReq) ! {
	if req.role_id == '' {
		return error('role_id is required')
	}
}

// ----------------- DTO 层 -----------------
pub struct DeleteTenantRoleReq {
	role_id string @[json: 'role_id']
}

pub struct DeleteTenantRoleResp {
	msg string @[json: 'msg']
}

// ----------------- Repository 层 -----------------
fn delete_role_repo(mut ctx Context, req DeleteTenantRoleReq) !DeleteTenantRoleResp {
	db, conn := ctx.dbpool.acquire() or { return error('Failed to acquire DB connection: ${err}') }
	defer {
		ctx.dbpool.release(conn) or { log.warn('Failed to release connection: ${err}') }
	}

	mut q := orm.new_query[CoreRole](db)
	q.set('del_flag = ?', 1)!.where('id = ?', req.role_id)!.update()!

	return DeleteTenantRoleResp{
		msg: 'Delete Tenant Role Successfully'
	}
}
