module db_api

pub const core_api = r"
REPLACE INTO `core_api` (`id`, `path`, `description`, `api_group`, `service_name`, `method`, `is_required`, `source_type`, `source_id`, `updater_id`, `updated_at`, `creator_id`, `created_at`, `del_flag`, `deleted_at`) VALUES
  ('00000000-0000-0000-0000-000000000001', '/core_api/admin/user/login', 'apiDesc.userLogin', 'user', 'Core', 'POST', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000002', '/core_api/admin/user/register', 'apiDesc.userRegister', 'user', 'Core', 'POST', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000003', '/core_api/admin/user/create', 'apiDesc.createUser', 'user', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000004', '/core_api/admin/user/update', 'apiDesc.updateUser', 'user', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000005', '/core_api/admin/user/change_password', 'apiDesc.userChangePassword', 'user', 'Core', 'POST', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000006', '/core_api/admin/user/info', 'apiDesc.userInfo', 'user', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000007', '/core_api/admin/user/list', 'apiDesc.userList', 'user', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000008', '/core_api/admin/user/delete', 'apiDesc.deleteUser', 'user', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000009', '/core_api/admin/user/perm', 'apiDesc.userPermissions', 'user', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000010', '/core_api/admin/user/profile', 'apiDesc.userProfile', 'user', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000011', '/core_api/admin/user/logout', 'apiDesc.logout', 'user', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000012', '/core_api/admin/user', 'apiDesc.getUserById', 'user', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000013', '/core_api/admin/user/refresh_token', 'apiDesc.refreshToken', 'user', 'Core', 'GET', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000014', '/core_api/admin/user/access_token', 'apiDesc.accessToken', 'user', 'Core', 'GET', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000015', '/core_api/admin/role/create', 'apiDesc.createRole', 'role', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000016', '/core_api/admin/role/update', 'apiDesc.updateRole', 'role', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000017', '/core_api/admin/role/delete', 'apiDesc.deleteRole', 'role', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000018', '/core_api/admin/role/list', 'apiDesc.roleList', 'role', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000019', '/core_api/admin/role', 'apiDesc.getRoleById', 'role', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000020', '/core_api/admin/menu/create', 'apiDesc.createMenu', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000021', '/core_api/admin/menu/update', 'apiDesc.updateMenu', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000022', '/core_api/admin/menu/delete', 'apiDesc.deleteMenu', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000023', '/core_api/admin/menu/list', 'apiDesc.menuList', 'menu', 'Core', 'GET', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000024', '/core_api/admin/menu/role/list', 'apiDesc.menuRoleList', 'authority', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000025', '/core_api/admin/menu_param/create', 'apiDesc.createMenuParam', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000026', '/core_api/admin/menu_param/update', 'apiDesc.updateMenuParam', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000027', '/core_api/admin/menu_param/list', 'apiDesc.menuParamListByMenuId', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000028', '/core_api/admin/menu_param/delete', 'apiDesc.deleteMenuParam', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000029', '/core_api/admin/menu_param', 'apiDesc.getMenuParamById', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000030', '/core_api/admin/menu', 'apiDesc.getMenuById', 'menu', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000031', '/core_api/admin/captcha', 'apiDesc.captcha', 'captcha', 'Core', 'GET', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000032', '/core_api/admin/authority/api/create_or_update', 'apiDesc.createOrUpdateApiAuthority', 'authority', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000033', '/core_api/admin/authority/api/role', 'apiDesc.APIAuthorityOfRole', 'authority', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000034', '/core_api/admin/authority/menu/create_or_update', 'apiDesc.createOrUpdateMenuAuthority', 'authority', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000035', '/core_api/admin/authority/menu/role', 'apiDesc.menuAuthorityOfRole', 'authority', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000036', '/core_api/admin/api/create', 'apiDesc.createApi', 'api', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000037', '/core_api/admin/api/update', 'apiDesc.updateApi', 'api', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000038', '/core_api/admin/api/delete', 'apiDesc.deleteAPI', 'api', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000039', '/core_api/admin/api/list', 'apiDesc.APIList', 'api', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000040', '/core_api/admin/api', 'apiDesc.getApiById', 'api', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000041', '/core_api/admin/oauth_provider/create', 'apiDesc.createProvider', 'oauth', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000042', '/core_api/admin/oauth_provider/update', 'apiDesc.updateProvider', 'oauth', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000043', '/core_api/admin/oauth_provider/delete', 'apiDesc.deleteProvider', 'oauth', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000044', '/core_api/admin/oauth_provider/list', 'apiDesc.getProviderList', 'oauth', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000045', '/core_api/admin/oauth/login', 'apiDesc.oauthLogin', 'oauth', 'Core', 'POST', 1, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000046', '/core_api/admin/oauth_provider', 'apiDesc.getProviderById', 'oauth', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000047', '/core_api/admin/token/create', 'apiDesc.createToken', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000048', '/core_api/admin/token/update', 'apiDesc.updateToken', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000049', '/core_api/admin/token/delete', 'apiDesc.deleteToken', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000050', '/core_api/admin/token/list', 'apiDesc.getTokenList', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000051', '/core_api/admin/token/logout', 'apiDesc.forceLoggingOut', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
  ('00000000-0000-0000-0000-000000000052', '/core_api/admin/token', 'apiDesc.getTokenById', 'token', 'Core', 'POST', 0, 'tenant', '00000000-0000-0000-0000-000000000000', NULL, '2024-11-18 00:54:02', NULL, '2024-11-18 00:54:02', 0, NULL);
"

pub const core_app = r'
'

pub const core_app_client = r'
'

pub const core_menu = r'
'

pub const core_project = r'
'

pub const core_role = r'
'

pub const core_role_api = r'
'

pub const core_role_menu = r'
'

pub const core_role_tenant_member = r'
'

pub const core_tenant = r'
'

pub const core_tenant_member = r'
'

pub const core_tenant_subapp = r'
'

pub const core_token = r'
'

pub const core_user = r'
'
